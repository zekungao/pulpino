
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00001D17,
    32'h844D0D13,
    32'h00001D97,
    32'h83CD8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h0C6000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'hCC221101,
    32'hCA266441,
    32'h147DCE06,
    32'h00EF4485,
    32'h8D6143A0,
    32'hFE951DE3,
    32'h46014681,
    32'h051345A1,
    32'h00EF09F0,
    32'h456136A0,
    32'h3B8000EF,
    32'h45014581,
    32'h394000EF,
    32'h45014581,
    32'h3E0000EF,
    32'h45E10068,
    32'h424000EF,
    32'h453240F2,
    32'h44D24462,
    32'h80826105,
    32'hCC221101,
    32'hCA266441,
    32'hC64EC84A,
    32'hCE06C452,
    32'h89AE8A2A,
    32'h147D8932,
    32'h00EF4485,
    32'h8D613DE0,
    32'hFE951DE3,
    32'h008A1613,
    32'h141346E1,
    32'h45A10059,
    32'h00EF450D,
    32'h852230A0,
    32'h358000EF,
    32'h45014581,
    32'h334000EF,
    32'h45014581,
    32'h380000EF,
    32'h854E85A2,
    32'h446240F2,
    32'h494244D2,
    32'h4A2249B2,
    32'h006F6105,
    32'h71593B60,
    32'hD6864505,
    32'hD2A6D4A2,
    32'hCECED0CA,
    32'hCAD6CCD2,
    32'hC6DEC8DA,
    32'hC2E6C4E2,
    32'hDE6EC0EA,
    32'h208000EF,
    32'h45014585,
    32'h40C000EF,
    32'h87936785,
    32'h0001BB87,
    32'hFFF517FD,
    32'h1A1027B7,
    32'hC3D84711,
    32'hF11FF0EF,
    32'h75138141,
    32'h07930FF5,
    32'h0B630EF0,
    32'h853700F5,
    32'h05930000,
    32'h05130230,
    32'h00EF7785,
    32'hA0014260,
    32'h00008537,
    32'h051345C5,
    32'h00EF79C5,
    32'h00EF4160,
    32'h46214660,
    32'h4501080C,
    32'hF25FF0EF,
    32'h4CF25782,
    32'h00008537,
    32'h5792C43E,
    32'h051345D5,
    32'hC63E7B05,
    32'h4AD249C2,
    32'h00EF5C32,
    32'h00EF3EA0,
    32'h596343A0,
    32'h69210990,
    32'h4A0164C1,
    32'h413A8AB3,
    32'h00008BB7,
    32'h7C890913,
    32'h00008B37,
    32'h440514FD,
    32'h8DB36D05,
    32'h00EF013A,
    32'h8D652D20,
    32'hFE851DE3,
    32'h00899613,
    32'h45A146E1,
    32'h00EF450D,
    32'h65212020,
    32'h250000EF,
    32'h45014581,
    32'h22C000EF,
    32'h45014581,
    32'h278000EF,
    32'h856E65A1,
    32'h2BC000EF,
    32'h85134599,
    32'h00EF734B,
    32'h55133820,
    32'h85A2004A,
    32'h00EF954A,
    32'h75133760,
    32'h85A200FA,
    32'h00EF954A,
    32'h0A0536A0,
    32'h05134599,
    32'h00EF73CB,
    32'h99EA35E0,
    32'h3AC000EF,
    32'hF94C99E3,
    32'h00008537,
    32'h051345B5,
    32'h00EF7445,
    32'h00EF3460,
    32'h5B633960,
    32'h49A20980,
    32'h692147B2,
    32'h4A0164C1,
    32'h00008BB7,
    32'h7C890913,
    32'h00008B37,
    32'h41378CB3,
    32'h440514FD,
    32'h8D336A85,
    32'h00EF013C,
    32'h8D6522A0,
    32'hFE851DE3,
    32'h00899613,
    32'h45A146E1,
    32'h00EF450D,
    32'h652115A0,
    32'h1A8000EF,
    32'h45014581,
    32'h184000EF,
    32'h45014581,
    32'h1D0000EF,
    32'h856A65A1,
    32'h214000EF,
    32'h85134599,
    32'h00EF734B,
    32'h55132DA0,
    32'h85A2004A,
    32'h00EF954A,
    32'h75132CE0,
    32'h85A200FA,
    32'h00EF954A,
    32'h0A052C20,
    32'h05134599,
    32'h00EF73CB,
    32'h99D62B60,
    32'h304000EF,
    32'hF94C19E3,
    32'h00008537,
    32'h02200593,
    32'h75450513,
    32'h29C000EF,
    32'h2EC000EF,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h50B60001,
    32'h54264501,
    32'h59065496,
    32'h4A6649F6,
    32'h4B464AD6,
    32'h4C264BB6,
    32'h4D064C96,
    32'h61655DF2,
    32'h00008082,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'h00912223,
    32'h2A8000EF,
    32'h00000593,
    32'h00E00513,
    32'h29C000EF,
    32'h00000593,
    32'h00D00513,
    32'h290000EF,
    32'h00000593,
    32'h00C00513,
    32'h284000EF,
    32'h04805E63,
    32'h00100493,
    32'h00000593,
    32'h01000513,
    32'h270000EF,
    32'h04940463,
    32'h00000593,
    32'h00B00513,
    32'h260000EF,
    32'h00200793,
    32'h02F40A63,
    32'h00000593,
    32'h00000513,
    32'h24C000EF,
    32'h00300793,
    32'h02F40063,
    32'h00048513,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h00000593,
    32'h01010113,
    32'h2280006F,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h01010113,
    32'h00008067,
    32'h00004737,
    32'hF0070713,
    32'h00869693,
    32'h02000793,
    32'h40B787B3,
    32'h00E6F6B3,
    32'h03F5F593,
    32'h1A102737,
    32'h00F51533,
    32'h00B6E5B3,
    32'h00A72423,
    32'h00C72623,
    32'h00B72823,
    32'h00008067,
    32'h01051513,
    32'h01059593,
    32'h01055513,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01072783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12783,
    32'h01051513,
    32'h01079793,
    32'h0107D793,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F72823,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00B795B3,
    32'h00A79533,
    32'h000017B7,
    32'hF0078793,
    32'h00F5F5B3,
    32'h0FF57513,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'h4055D793,
    32'hFF010113,
    32'h7FF7F793,
    32'h01F5F593,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12683,
    32'h00812783,
    32'h1A102737,
    32'h00070813,
    32'h04F6D063,
    32'h00072783,
    32'h4107D793,
    32'h0FF7F793,
    32'hFE078AE3,
    32'h00C12783,
    32'h02082583,
    32'h00C12683,
    32'h00279793,
    32'h00168693,
    32'h00D12623,
    32'h00C12603,
    32'h00812683,
    32'h00F507B3,
    32'h00B7A023,
    32'hFCD644E3,
    32'h01010113,
    32'h00008067,
    32'h1A1076B7,
    32'h0046A703,
    32'h1A1007B7,
    32'h00276713,
    32'h00E6A223,
    32'h08300713,
    32'h00E7A623,
    32'h0085D613,
    32'h0A700713,
    32'h0FF5F593,
    32'h00C7A223,
    32'h00B7A023,
    32'h00E7A423,
    32'h00300713,
    32'h00E7A623,
    32'h0047A703,
    32'h0F077713,
    32'h00276713,
    32'h00E7A223,
    32'h00008067,
    32'h04058863,
    32'h1A1006B7,
    32'h0146A783,
    32'h0207F793,
    32'hFE078CE3,
    32'h00054603,
    32'h1A100737,
    32'h00150793,
    32'h00C72023,
    32'hFFF58593,
    32'h04050513,
    32'h0140006F,
    32'hFFF7C703,
    32'hFFF58593,
    32'h00E6A023,
    32'h00A78863,
    32'h00178793,
    32'hFE0596E3,
    32'h00008067,
    32'hFA059EE3,
    32'h00008067,
    32'h1A100737,
    32'h01472783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00C12703,
    32'h00A797B3,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00A595B3,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F6A023,
    32'h00008067,
    32'h636F6C42,
    32'h0000206B,
    32'h6E6F6420,
    32'h00000A65,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h4F525245,
    32'h57203A52,
    32'h6F626E69,
    32'h5320646E,
    32'h66204950,
    32'h6873616C,
    32'h746F6E20,
    32'h756F6620,
    32'h000A646E,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h0000001C,
    32'h00000018,
    32'hFFFFF95C,
    32'h00000050,
    32'h200E4200,
    32'h7E081142,
    32'h7D091146,
    32'h007F0111,
    32'h00000024,
    32'h00000038,
    32'hFFFFF98C,
    32'h00000062,
    32'h200E4200,
    32'h7E081142,
    32'h7D09114C,
    32'h117C1211,
    32'h14117B13,
    32'h7F01117A,
    32'h00000038,
    32'h00000060,
    32'hFFFFF9C6,
    32'h00000224,
    32'h700E4200,
    32'h7F01115C,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h16117915,
    32'h77171178,
    32'h11761811,
    32'h1A117519,
    32'h731B1174,
    32'h0000001C,
    32'h0000009C,
    32'hFFFFFBB0,
    32'h000000B4,
    32'h100E4400,
    32'h7E081148,
    32'h7F011150,
    32'h007D0911};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule